class alu_driver extends uvm_driver#(alu_sequence_item);
  `uvm_component_utils(alu_driver);
  virtual alu_interface vif;
  alu_sequence_item item;
  function new(string name="alu_driver", uvm_component parent);
    super.new(name,parent);
  endfunction
  
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
       if(!(uvm_config_db #(virtual alu_interface)::get(this, "*", "vif", vif))) begin
      `uvm_error("DRIVER_CLASS", "Failed to get VIF from config DB!")
    end	
  endfunction:build_phase
  
  
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
 
  endfunction: connect_phase
  
  
  task run_phase(uvm_phase phase);
    super.run_phase(phase);
    
    
    forever begin
      item = alu_sequence_item::type_id::create("item");
      seq_item_port.get_next_item(item);
      
      drive(item);
      seq_item_port.item_done();
      
    end
  endtask: run_phase
  
  
  
  task drive(alu_sequence_item item);
    @(posedge vif.clock)
    	vif.reset<=item.reset;
    	vif.A<= item.A;
    	vif.B<=item.B;
    	vif.op <=item.op;
  endtask: drive
  
endclass:alu_driver;